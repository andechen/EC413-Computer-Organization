`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/13/2021 06:55:55 PM
// Design Name: 
// Module Name: NBitSLT
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module NBitSLT_str#(
    parameter N = 32
)(
    output [N-1:0] out,
    input  [N-1:0] input1,
    input  [N-1:0] input2
    );
    
    // if input1 < input 2, out is 1 else out is 0
    // 
    
endmodule
