`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/12/2021 05:52:59 PM
// Design Name: 
// Module Name: top_str
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top_str(
    input [N-1:0] a,
    input [N-1:0] b,
    input c_in,
    input [N-1:0] sum,
    input c_out
    );
    
    // mux that chooses between doing the NOT of a and adding a and b
    
endmodule
